LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity reg8b_serial IS
	

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TP1EX1 IS
	PORT (  E1, E0		: in STD_LOGIC;
		S3, S2, S1, S0	: OUT STD_LOGIC);
END ENTITY TP1EX1;

ARCHITECTURE fdd_TP1EX1 OF TP1EX1 IS
	SIGNAL S : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SUBTYPE selecteur IS STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
	(S3, S2 ,S1, S0) <= S;
	WITH selecteur'(E1 & E0) SELECT
		S <=	"0001" WHEN "00",
			"0010" WHEN "01",
			"0100" WHEN "10",
			"1000" WHEN "11",
			"0000" WHEN OTHERS;
END ARCHITECTURE fdd_TP1EX1;

--Ce code correspond à un décodeur 2->4
